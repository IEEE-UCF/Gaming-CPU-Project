module axi_dcache_port #(
  // TODO: Parameter setups
  parameter unsigned 
)(
  // TODO: Port set up
  ports

  // TODO: Input logic
  input logic clk_i,
  input logic rst_ni
  
  
);

endmodule

