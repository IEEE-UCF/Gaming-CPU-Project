module axi_icache_port #(
  // TODO: Parameter setups
  parameter
)(
  // TODO: Port set up
  ports

  // TODO: Input logic
  input logic clk_i,
  input logic rst_ni
  
);

endmodule
