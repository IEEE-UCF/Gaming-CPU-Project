module cache_miss_unit #(
    parameters
) (
    ports
);

endmodule
