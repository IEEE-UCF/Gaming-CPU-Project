module cache_tags #(
    parameters
) (
    ports
);

endmodule
