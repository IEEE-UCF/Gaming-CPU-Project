//Divyesh Narra