module axi_dcache_port #(
  parameter
)(
  ports
);

endmodule
