module cache_coherency_none #(
    parameters
) (
    ports
);

endmodule