module axi_to_axi_lite #(
  // TODO: Parameter setups
  parameter
)(
  // TODO: Port set up
  ports

  // TODO: Input logic
  input logic clk_i,
  input logic rst_ni
  
);

endmodule
