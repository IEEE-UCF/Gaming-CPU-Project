/***************************RECEIVE rx_i*******************************/
// Serial input -> shift register -> FIFO

/***************************FIFO MANAGEMENT****************************/
// Push/pop data, update pointers and count
