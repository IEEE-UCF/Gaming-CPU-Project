module dcache #(
    parameter int INSTR_WIDTH = 32,
    parameter ADDR_WIDTH = 32,
    parameter LINE_SIZE = 64,
    parameter WAYS = 4,
    parameter DMEM_SIZE = 16384
) (
    ports
);

endmodule