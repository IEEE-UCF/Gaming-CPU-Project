//Divyesh