module l2_cache #(
    parameter int INSTR_WIDTH = 32,
    parameter int ADDR_WIDTH = 32,
    parameter int LINE_SIZE = 64,
    parameter int WAYS = 4,
    parameter int L2_SIZE = 262144
) (
    ports
);

endmodule