//
//
//

package interconnect_pkg;
  
  parameter int unsigned ADDR_WIDTH = 32;
  parameter int unsigned DATA_WIDTH = 64;
  
endpackage
