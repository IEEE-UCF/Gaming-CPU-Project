/***************************RECEIVE rx_i*******************************/
// Serial input -> shift register -> FIFO
