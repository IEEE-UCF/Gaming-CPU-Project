//


package interconnect_pkg;

// AXI Data Widths
parameter int unsigned AXI_ADDR_WIDTH = 32;
parameter int unsigned AXI_DATA_WIDTH = 64;
parameter int unsigned AXI_ID_WIDTH = 4;
parameter int unsigned AXI_USER_WIDTH = 1;

parameter int unsigned AXI_STRB_WIDTH = AXI_DATA_WIDTH/8;

// Master IDs (TBD)

// Address Map (TBD)

// Cache Line

    
endpackage